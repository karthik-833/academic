module fifo #(
    parameter DATA_WIDTH = 8,  // Data bus width  
    parameter DEPTH = 16       // FIFO depth (number of entries)  
)(
    input  logic                     clk,       // Clock signal  
    input  logic                     rst,       // Synchronous reset (active high)  
    input  logic                     wr_en,     // Write enable signal  
    input  logic                     rd_en,     // Read enable signal  
    input  logic [DATA_WIDTH-1:0]    data_in,   // Input data  
    output logic [DATA_WIDTH-1:0]    data_out,  // Output data  
    output logic                     empty,     // FIFO is empty  
    output logic                     full    );   // FIFO is full);

    // Internal storage and pointers
    logic [DATA_WIDTH-1:0] mem[0:DEPTH-1]; // Memory array
    logic [$clog2(DEPTH)-1:0] wr_ptr, rd_ptr,pr ,pw; // Write and read pointers
    logic [$clog2(DEPTH)-1:0] count;   
    logic write;
    logic read;
    // Tracks the number of entries in the FIFO
    assign full  = (count == DEPTH);
    assign empty = (count == 0);
    assign read = (rd_en && !empty);
    assign write = (wr_en && !full && (!(rd_ptr == wr_ptr) || read));
    

    // Write logic
    always_ff @(posedge clk) begin
          wr_ptr = pw;
        if (rst) begin
            wr_ptr = 0;
        end else if (write) begin
          mem[wr_ptr] = data_in;
            pw = wr_ptr + 1;
        end
    end

    // Read logic
    always_ff @(posedge clk) begin
        rd_ptr=pr;
        if (rst) begin
            rd_ptr = 0;
  end else if (read)  begin
           data_out = mem[rd_ptr];
            pr = rd_ptr + 1;
        end
    end

    // Count tracking
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            count = 0;
        end else if (wr_en && !full && rd_en && !empty) begin
            count <= count; // Simultaneous read and write
        end else if (wr_en && !full) begin
            count = count + 1;
        end else if (rd_en && !empty) begin
            count = count - 1;
        end
    end

  // Ensure data is written only when FIFO is not full
always @(posedge clk) begin
    if (rst) begin
        assert property (1);  // No violations during reset
    end else begin
        assert property (write ? ((!wr_en) || (!full)) : 1'b1); // Write occurs only if FIFO is not full
    end
end

// Ensure data is read only when FIFO is not empty
always @(posedge clk) begin
    if (rst) begin
        assert property (1);  // No violations during reset
    end else begin
        assert property (read ? (!(empty && rd_en)): 1'b1);  // Read occurs only if FIFO is not empty
    end
end

// Count must always be between 0 and DEPTH
always @(posedge clk) begin
    if (rst) begin
        assert property (count == 0); // Ensure count is reset to 0
    end else begin
        assert property (count >= 0 && count <= DEPTH);  // Assert count is in valid range
    end
end

// Data integrity check for matching written and read data
always @(posedge clk) begin
    if (rst) begin
        assert property (1); // No violations during reset
    end else begin
       // assert property ((rd_ptr ==  wr_ptr) ? ((rd_en && wr_en ) ? (data_in == data_out): 1'b1)  : 1'b1) ; // Write and read match on the same cycle
    end
end

// No writing occurs when FIFO is full
always @(posedge clk) begin
    if (rst) begin
        assert property (1);  // No violations during reset
    end else begin
        assert property (!(full && wr_en)); // No write when FIFO is full
    end
end
// Ensure new data is not written until the old data is read
always @(posedge clk) begin
    if (rst) begin
        assert property (1); // No violations during reset
    end else begin
        // If the FIFO is not empty, write should not overtake read
        assert property (!(write && (wr_ptr == rd_ptr) && !read)); 
    end
end



endmodule
